�      �   �     "�   �     H�   �     e�   �     l�   �     l�   �     o�   �      �   �     W�   �     o�   �     r�   �     l�   �     d�   �     "�   